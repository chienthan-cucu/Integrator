module add_signed_5_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A;
  input [21:0] B;
  output [21:0] Z;
  wire [20:0] A;
  wire [21:0] B;
  wire [21:0] Z;
  wire n_69, n_72, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_179;
  nand g4 (n_72, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_69, B[9], n_116);
  nand g61 (n_120, n_117, n_118, n_69);
  xor g62 (n_119, A[9], B[9]);
  xor g63 (Z[9], n_116, n_119);
  nand g64 (n_121, A[10], B[10]);
  nand g65 (n_122, A[10], n_120);
  nand g66 (n_123, B[10], n_120);
  nand g67 (n_125, n_121, n_122, n_123);
  xor g68 (n_124, A[10], B[10]);
  xor g69 (Z[10], n_120, n_124);
  nand g70 (n_126, A[11], B[11]);
  nand g71 (n_127, A[11], n_125);
  nand g72 (n_128, B[11], n_125);
  nand g73 (n_130, n_126, n_127, n_128);
  xor g74 (n_129, A[11], B[11]);
  xor g75 (Z[11], n_125, n_129);
  nand g76 (n_131, A[12], B[12]);
  nand g77 (n_132, A[12], n_130);
  nand g78 (n_133, B[12], n_130);
  nand g79 (n_135, n_131, n_132, n_133);
  xor g80 (n_134, A[12], B[12]);
  xor g81 (Z[12], n_130, n_134);
  nand g82 (n_136, A[13], B[13]);
  nand g83 (n_137, A[13], n_135);
  nand g84 (n_138, B[13], n_135);
  nand g85 (n_140, n_136, n_137, n_138);
  xor g86 (n_139, A[13], B[13]);
  xor g87 (Z[13], n_135, n_139);
  nand g88 (n_141, A[14], B[14]);
  nand g89 (n_142, A[14], n_140);
  nand g90 (n_143, B[14], n_140);
  nand g91 (n_145, n_141, n_142, n_143);
  xor g92 (n_144, A[14], B[14]);
  xor g93 (Z[14], n_140, n_144);
  nand g94 (n_146, A[15], B[15]);
  nand g95 (n_147, A[15], n_145);
  nand g96 (n_148, B[15], n_145);
  nand g97 (n_150, n_146, n_147, n_148);
  xor g98 (n_149, A[15], B[15]);
  xor g99 (Z[15], n_145, n_149);
  nand g100 (n_151, A[16], B[16]);
  nand g101 (n_152, A[16], n_150);
  nand g102 (n_153, B[16], n_150);
  nand g103 (n_155, n_151, n_152, n_153);
  xor g104 (n_154, A[16], B[16]);
  xor g105 (Z[16], n_150, n_154);
  nand g106 (n_156, A[17], B[17]);
  nand g107 (n_157, A[17], n_155);
  nand g108 (n_158, B[17], n_155);
  nand g109 (n_160, n_156, n_157, n_158);
  xor g110 (n_159, A[17], B[17]);
  xor g111 (Z[17], n_155, n_159);
  nand g112 (n_161, A[18], B[18]);
  nand g113 (n_162, A[18], n_160);
  nand g114 (n_163, B[18], n_160);
  nand g115 (n_165, n_161, n_162, n_163);
  xor g116 (n_164, A[18], B[18]);
  xor g117 (Z[18], n_160, n_164);
  nand g118 (n_166, A[19], B[19]);
  nand g119 (n_167, A[19], n_165);
  nand g120 (n_168, B[19], n_165);
  nand g121 (n_170, n_166, n_167, n_168);
  xor g122 (n_169, A[19], B[19]);
  xor g123 (Z[19], n_165, n_169);
  nand g124 (n_171, A[20], B[20]);
  nand g125 (n_172, A[20], n_170);
  nand g126 (n_173, B[20], n_170);
  nand g127 (n_175, n_171, n_172, n_173);
  xor g128 (n_174, A[20], B[20]);
  xor g129 (Z[20], n_170, n_174);
  xor g135 (Z[21], n_175, n_179);
  xor g137 (n_179, A[20], B[21]);
  or g138 (n_78, wc, n_72);
  not gc (wc, A[1]);
  or g139 (n_79, wc0, n_72);
  not gc0 (wc0, B[1]);
  xnor g140 (Z[1], n_72, n_80);
endmodule

module add_signed_5_GENERIC(A, B, Z);
  input [20:0] A;
  input [21:0] B;
  output [21:0] Z;
  wire [20:0] A;
  wire [21:0] B;
  wire [21:0] Z;
  add_signed_5_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module csa_tree_add_125_31_group_301_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( ( 367 * $signed(in_1) )  + ( 1314 * $signed(in_2) )  )  + ( 367 * $signed(in_0) )  )  ;"
  input [20:0] in_0;
  input [21:0] in_1, in_2;
  output [20:0] out_0;
  wire [20:0] in_0;
  wire [21:0] in_1, in_2;
  wire [20:0] out_0;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_138, n_143;
  wire n_144, n_145, n_149, n_150, n_151, n_152, n_153, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_410;
  wire n_411, n_412, n_413, n_414, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_454, n_455, n_456, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_928, n_933, n_938;
  wire n_943, n_948, n_953, n_958, n_963, n_968, n_973, n_981;
  wire n_983, n_986, n_987, n_988, n_989, n_990, n_991, n_993;
  wire n_994, n_995, n_996, n_997, n_999, n_1000, n_1001, n_1002;
  wire n_1003, n_1005, n_1006, n_1007, n_1008, n_1009, n_1011, n_1012;
  wire n_1013, n_1014, n_1015, n_1017, n_1018, n_1019, n_1020, n_1021;
  wire n_1023, n_1024, n_1025, n_1026, n_1027, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1035, n_1036, n_1037, n_1038, n_1039, n_1041;
  wire n_1042, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1051;
  wire n_1053, n_1055, n_1056, n_1058, n_1059, n_1061, n_1063, n_1065;
  wire n_1066, n_1068, n_1069, n_1071, n_1073, n_1075, n_1076, n_1078;
  wire n_1079, n_1081, n_1083, n_1085, n_1086, n_1088, n_1090, n_1091;
  wire n_1092, n_1094, n_1095, n_1096, n_1098, n_1099, n_1100, n_1101;
  wire n_1103, n_1105, n_1107, n_1108, n_1109, n_1111, n_1112, n_1113;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1121, n_1122, n_1123;
  wire n_1125, n_1126, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133;
  wire n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141;
  wire n_1143, n_1144, n_1145, n_1147, n_1148, n_1150, n_1151, n_1152;
  wire n_1154, n_1155, n_1156, n_1158, n_1159, n_1160, n_1161, n_1163;
  wire n_1164, n_1165, n_1167, n_1168, n_1169, n_1170, n_1172, n_1173;
  wire n_1175, n_1176, n_1178, n_1179, n_1180, n_1181, n_1183, n_1184;
  wire n_1185, n_1187, n_1188, n_1189, n_1190, n_1192, n_1193, n_1195;
  wire n_1196;
  nand g196 (n_104, n_412, n_413, n_414);
  nand g202 (n_138, n_416, n_417, n_418);
  nand g208 (n_143, n_420, n_421, n_422);
  xor g210 (n_124, n_423, n_138);
  nand g214 (n_102, n_424, n_425, n_426);
  nand g222 (n_149, n_428, n_429, n_430);
  xor g224 (n_145, n_431, in_0[5]);
  nand g227 (n_434, in_2[0], in_0[5]);
  nand g228 (n_152, n_410, n_433, n_434);
  xor g229 (n_435, n_143, n_144);
  xor g230 (n_123, n_435, n_145);
  nand g231 (n_436, n_143, n_144);
  nand g232 (n_437, n_145, n_144);
  nand g233 (n_438, n_143, n_145);
  nand g234 (n_101, n_436, n_437, n_438);
  nand g240 (n_157, n_440, n_441, n_442);
  nand g246 (n_156, n_444, n_414, n_446);
  xor g248 (n_153, n_447, n_150);
  nand g250 (n_449, n_150, n_149);
  nand g252 (n_161, n_448, n_449, n_450);
  xor g253 (n_451, n_151, n_152);
  xor g254 (n_122, n_451, n_153);
  nand g255 (n_452, n_151, n_152);
  nand g256 (n_453, n_153, n_152);
  nand g257 (n_454, n_151, n_153);
  nand g258 (n_100, n_452, n_453, n_454);
  nand g264 (n_166, n_456, n_416, n_458);
  xor g266 (n_159, n_459, in_1[0]);
  nand g270 (n_165, n_460, n_461, n_462);
  xor g271 (n_463, in_2[6], in_0[0]);
  xor g272 (n_160, n_463, n_156);
  nand g273 (n_464, in_2[6], in_0[0]);
  nand g274 (n_465, n_156, in_0[0]);
  nand g275 (n_466, in_2[6], n_156);
  nand g276 (n_170, n_464, n_465, n_466);
  xor g277 (n_467, n_157, n_158);
  xor g278 (n_162, n_467, n_159);
  nand g279 (n_468, n_157, n_158);
  nand g280 (n_469, n_159, n_158);
  nand g281 (n_470, n_157, n_159);
  nand g282 (n_172, n_468, n_469, n_470);
  xor g283 (n_471, n_160, n_161);
  xor g284 (n_121, n_471, n_162);
  nand g285 (n_472, n_160, n_161);
  nand g286 (n_473, n_162, n_161);
  nand g287 (n_474, n_160, n_162);
  nand g288 (n_99, n_472, n_473, n_474);
  nand g294 (n_179, n_476, n_477, n_478);
  xor g296 (n_169, n_419, in_0[0]);
  nand g298 (n_481, in_0[0], in_2[3]);
  nand g300 (n_178, n_420, n_481, n_482);
  xor g302 (n_167, n_483, in_2[7]);
  nand g305 (n_486, in_1[1], in_2[7]);
  nand g306 (n_177, n_484, n_485, n_486);
  xor g307 (n_487, in_1[0], in_0[1]);
  xor g308 (n_171, n_487, n_165);
  nand g309 (n_488, in_1[0], in_0[1]);
  nand g310 (n_489, n_165, in_0[1]);
  nand g311 (n_490, in_1[0], n_165);
  nand g312 (n_183, n_488, n_489, n_490);
  xor g313 (n_491, n_166, n_167);
  xor g314 (n_173, n_491, n_168);
  nand g315 (n_492, n_166, n_167);
  nand g316 (n_493, n_168, n_167);
  nand g317 (n_494, n_166, n_168);
  nand g318 (n_185, n_492, n_493, n_494);
  xor g319 (n_495, n_169, n_170);
  xor g320 (n_174, n_495, n_171);
  nand g321 (n_496, n_169, n_170);
  nand g322 (n_497, n_171, n_170);
  nand g323 (n_498, n_169, n_171);
  nand g324 (n_188, n_496, n_497, n_498);
  xor g325 (n_499, n_172, n_173);
  xor g326 (n_120, n_499, n_174);
  nand g327 (n_500, n_172, n_173);
  nand g328 (n_501, n_174, n_173);
  nand g329 (n_502, n_172, n_174);
  nand g330 (n_98, n_500, n_501, n_502);
  nand g336 (n_192, n_504, n_505, n_506);
  nand g340 (n_509, in_0[1], in_2[4]);
  nand g342 (n_193, n_508, n_509, n_510);
  xor g344 (n_182, n_511, in_2[8]);
  nand g347 (n_514, in_1[2], in_2[8]);
  nand g348 (n_194, n_512, n_513, n_514);
  xor g349 (n_515, in_1[1], in_0[2]);
  xor g350 (n_184, n_515, n_177);
  nand g351 (n_516, in_1[1], in_0[2]);
  nand g352 (n_517, n_177, in_0[2]);
  nand g353 (n_518, in_1[1], n_177);
  nand g354 (n_199, n_516, n_517, n_518);
  xor g355 (n_519, n_178, n_179);
  xor g356 (n_186, n_519, n_180);
  nand g357 (n_520, n_178, n_179);
  nand g358 (n_521, n_180, n_179);
  nand g359 (n_522, n_178, n_180);
  nand g360 (n_200, n_520, n_521, n_522);
  xor g361 (n_523, n_181, n_182);
  xor g362 (n_187, n_523, n_183);
  nand g363 (n_524, n_181, n_182);
  nand g364 (n_525, n_183, n_182);
  nand g365 (n_526, n_181, n_183);
  nand g366 (n_203, n_524, n_525, n_526);
  xor g367 (n_527, n_184, n_185);
  xor g368 (n_189, n_527, n_186);
  nand g369 (n_528, n_184, n_185);
  nand g370 (n_529, n_186, n_185);
  nand g371 (n_530, n_184, n_186);
  nand g372 (n_204, n_528, n_529, n_530);
  xor g373 (n_531, n_187, n_188);
  xor g374 (n_119, n_531, n_189);
  nand g375 (n_532, n_187, n_188);
  nand g376 (n_533, n_189, n_188);
  nand g377 (n_534, n_187, n_189);
  nand g378 (n_97, n_532, n_533, n_534);
  nand g384 (n_213, n_536, n_537, n_538);
  xor g385 (n_539, in_0[3], in_2[2]);
  nand g387 (n_540, in_0[3], in_2[2]);
  nand g390 (n_210, n_540, n_541, n_542);
  xor g392 (n_198, n_543, in_2[5]);
  nand g395 (n_546, in_1[2], in_2[5]);
  nand g396 (n_212, n_544, n_545, n_546);
  xor g397 (n_547, in_2[9], in_1[3]);
  xor g398 (n_197, n_547, in_0[2]);
  nand g399 (n_548, in_2[9], in_1[3]);
  nand g400 (n_549, in_0[2], in_1[3]);
  nand g401 (n_550, in_2[9], in_0[2]);
  nand g402 (n_211, n_548, n_549, n_550);
  xor g403 (n_551, n_192, n_193);
  xor g404 (n_201, n_551, n_194);
  nand g405 (n_552, n_192, n_193);
  nand g406 (n_553, n_194, n_193);
  nand g407 (n_554, n_192, n_194);
  nand g408 (n_217, n_552, n_553, n_554);
  xor g409 (n_555, n_195, n_196);
  xor g410 (n_202, n_555, n_197);
  nand g411 (n_556, n_195, n_196);
  nand g412 (n_557, n_197, n_196);
  nand g413 (n_558, n_195, n_197);
  nand g414 (n_220, n_556, n_557, n_558);
  xor g415 (n_559, n_198, n_199);
  xor g416 (n_205, n_559, n_200);
  nand g417 (n_560, n_198, n_199);
  nand g418 (n_561, n_200, n_199);
  nand g419 (n_562, n_198, n_200);
  nand g420 (n_223, n_560, n_561, n_562);
  xor g421 (n_563, n_201, n_202);
  xor g422 (n_206, n_563, n_203);
  nand g423 (n_564, n_201, n_202);
  nand g424 (n_565, n_203, n_202);
  nand g425 (n_566, n_201, n_203);
  nand g426 (n_224, n_564, n_565, n_566);
  xor g427 (n_567, n_204, n_205);
  xor g428 (n_118, n_567, n_206);
  nand g429 (n_568, n_204, n_205);
  nand g430 (n_569, n_206, n_205);
  nand g431 (n_570, n_204, n_206);
  nand g432 (n_96, n_568, n_569, n_570);
  xor g436 (n_216, n_571, in_2[3]);
  nand g438 (n_573, in_2[3], in_0[4]);
  nand g440 (n_229, n_572, n_573, n_574);
  nand g446 (n_230, n_576, n_577, n_578);
  xor g447 (n_579, in_2[6], in_2[10]);
  xor g448 (n_214, n_579, in_1[4]);
  nand g449 (n_580, in_2[6], in_2[10]);
  nand g450 (n_581, in_1[4], in_2[10]);
  nand g451 (n_582, in_2[6], in_1[4]);
  nand g452 (n_231, n_580, n_581, n_582);
  xor g453 (n_583, in_0[3], n_209);
  xor g454 (n_218, n_583, n_210);
  nand g455 (n_584, in_0[3], n_209);
  nand g456 (n_585, n_210, n_209);
  nand g457 (n_586, in_0[3], n_210);
  nand g458 (n_237, n_584, n_585, n_586);
  xor g459 (n_587, n_211, n_212);
  xor g460 (n_219, n_587, n_213);
  nand g461 (n_588, n_211, n_212);
  nand g462 (n_589, n_213, n_212);
  nand g463 (n_590, n_211, n_213);
  nand g464 (n_236, n_588, n_589, n_590);
  xor g465 (n_591, n_214, n_215);
  xor g466 (n_221, n_591, n_216);
  nand g467 (n_592, n_214, n_215);
  nand g468 (n_593, n_216, n_215);
  nand g469 (n_594, n_214, n_216);
  nand g470 (n_238, n_592, n_593, n_594);
  xor g471 (n_595, n_217, n_218);
  xor g472 (n_222, n_595, n_219);
  nand g473 (n_596, n_217, n_218);
  nand g474 (n_597, n_219, n_218);
  nand g475 (n_598, n_217, n_219);
  nand g476 (n_242, n_596, n_597, n_598);
  xor g477 (n_599, n_220, n_221);
  xor g478 (n_225, n_599, n_222);
  nand g479 (n_600, n_220, n_221);
  nand g480 (n_601, n_222, n_221);
  nand g481 (n_602, n_220, n_222);
  nand g482 (n_245, n_600, n_601, n_602);
  xor g483 (n_603, n_223, n_224);
  xor g484 (n_117, n_603, n_225);
  nand g485 (n_604, n_223, n_224);
  nand g486 (n_605, n_225, n_224);
  nand g487 (n_606, n_223, n_225);
  nand g488 (n_95, n_604, n_605, n_606);
  nand g494 (n_248, n_608, n_609, n_610);
  xor g495 (n_611, in_0[5], in_2[4]);
  nand g497 (n_612, in_0[5], in_2[4]);
  nand g500 (n_249, n_612, n_613, n_614);
  xor g502 (n_234, n_615, in_2[7]);
  nand g505 (n_618, in_1[4], in_2[7]);
  nand g506 (n_251, n_616, n_617, n_618);
  xor g507 (n_619, in_2[11], in_1[5]);
  xor g508 (n_232, n_619, in_0[4]);
  nand g509 (n_620, in_2[11], in_1[5]);
  nand g510 (n_621, in_0[4], in_1[5]);
  nand g511 (n_622, in_2[11], in_0[4]);
  nand g512 (n_250, n_620, n_621, n_622);
  xor g513 (n_623, n_228, n_229);
  xor g514 (n_239, n_623, n_230);
  nand g515 (n_624, n_228, n_229);
  nand g516 (n_625, n_230, n_229);
  nand g517 (n_626, n_228, n_230);
  nand g518 (n_256, n_624, n_625, n_626);
  xor g519 (n_627, n_231, n_232);
  xor g520 (n_240, n_627, n_233);
  nand g521 (n_628, n_231, n_232);
  nand g522 (n_629, n_233, n_232);
  nand g523 (n_630, n_231, n_233);
  nand g524 (n_257, n_628, n_629, n_630);
  xor g525 (n_631, n_234, n_235);
  xor g526 (n_241, n_631, n_236);
  nand g527 (n_632, n_234, n_235);
  nand g528 (n_633, n_236, n_235);
  nand g529 (n_634, n_234, n_236);
  nand g530 (n_261, n_632, n_633, n_634);
  xor g531 (n_635, n_237, n_238);
  xor g532 (n_243, n_635, n_239);
  nand g533 (n_636, n_237, n_238);
  nand g534 (n_637, n_239, n_238);
  nand g535 (n_638, n_237, n_239);
  nand g536 (n_262, n_636, n_637, n_638);
  xor g537 (n_639, n_240, n_241);
  xor g538 (n_244, n_639, n_242);
  nand g539 (n_640, n_240, n_241);
  nand g540 (n_641, n_242, n_241);
  nand g541 (n_642, n_240, n_242);
  nand g542 (n_265, n_640, n_641, n_642);
  xor g543 (n_643, n_243, n_244);
  xor g544 (n_116, n_643, n_245);
  nand g545 (n_644, n_243, n_244);
  nand g546 (n_645, n_245, n_244);
  nand g547 (n_646, n_243, n_245);
  nand g548 (n_94, n_644, n_645, n_646);
  nand g554 (n_268, n_648, n_649, n_650);
  xor g555 (n_651, in_0[6], in_2[5]);
  nand g557 (n_652, in_0[6], in_2[5]);
  nand g560 (n_269, n_652, n_653, n_654);
  xor g562 (n_253, n_655, in_2[8]);
  nand g565 (n_658, in_1[5], in_2[8]);
  nand g566 (n_271, n_656, n_657, n_658);
  xor g567 (n_659, in_2[12], in_1[6]);
  xor g568 (n_255, n_659, in_0[5]);
  nand g569 (n_660, in_2[12], in_1[6]);
  nand g570 (n_661, in_0[5], in_1[6]);
  nand g571 (n_662, in_2[12], in_0[5]);
  nand g572 (n_270, n_660, n_661, n_662);
  xor g573 (n_663, n_248, n_249);
  xor g574 (n_258, n_663, n_250);
  nand g575 (n_664, n_248, n_249);
  nand g576 (n_665, n_250, n_249);
  nand g577 (n_666, n_248, n_250);
  nand g578 (n_276, n_664, n_665, n_666);
  xor g579 (n_667, n_251, n_252);
  xor g580 (n_259, n_667, n_253);
  nand g581 (n_668, n_251, n_252);
  nand g582 (n_669, n_253, n_252);
  nand g583 (n_670, n_251, n_253);
  nand g584 (n_277, n_668, n_669, n_670);
  xor g585 (n_671, n_254, n_255);
  xor g586 (n_260, n_671, n_256);
  nand g587 (n_672, n_254, n_255);
  nand g588 (n_673, n_256, n_255);
  nand g589 (n_674, n_254, n_256);
  nand g590 (n_281, n_672, n_673, n_674);
  xor g591 (n_675, n_257, n_258);
  xor g592 (n_263, n_675, n_259);
  nand g593 (n_676, n_257, n_258);
  nand g594 (n_677, n_259, n_258);
  nand g595 (n_678, n_257, n_259);
  nand g596 (n_282, n_676, n_677, n_678);
  xor g597 (n_679, n_260, n_261);
  xor g598 (n_264, n_679, n_262);
  nand g599 (n_680, n_260, n_261);
  nand g600 (n_681, n_262, n_261);
  nand g601 (n_682, n_260, n_262);
  nand g602 (n_284, n_680, n_681, n_682);
  xor g603 (n_683, n_263, n_264);
  xor g604 (n_115, n_683, n_265);
  nand g605 (n_684, n_263, n_264);
  nand g606 (n_685, n_265, n_264);
  nand g607 (n_686, n_263, n_265);
  nand g608 (n_93, n_684, n_685, n_686);
  nand g614 (n_288, n_688, n_689, n_690);
  xor g615 (n_691, in_0[7], in_2[6]);
  nand g617 (n_692, in_0[7], in_2[6]);
  nand g620 (n_289, n_692, n_693, n_694);
  xor g622 (n_273, n_695, in_2[9]);
  nand g625 (n_698, in_1[6], in_2[9]);
  nand g626 (n_291, n_696, n_697, n_698);
  xor g627 (n_699, in_2[13], in_1[7]);
  xor g628 (n_275, n_699, in_0[6]);
  nand g629 (n_700, in_2[13], in_1[7]);
  nand g630 (n_701, in_0[6], in_1[7]);
  nand g631 (n_702, in_2[13], in_0[6]);
  nand g632 (n_290, n_700, n_701, n_702);
  xor g633 (n_703, n_268, n_269);
  xor g634 (n_278, n_703, n_270);
  nand g635 (n_704, n_268, n_269);
  nand g636 (n_705, n_270, n_269);
  nand g637 (n_706, n_268, n_270);
  nand g638 (n_296, n_704, n_705, n_706);
  xor g639 (n_707, n_271, n_272);
  xor g640 (n_279, n_707, n_273);
  nand g641 (n_708, n_271, n_272);
  nand g642 (n_709, n_273, n_272);
  nand g643 (n_710, n_271, n_273);
  nand g644 (n_297, n_708, n_709, n_710);
  xor g645 (n_711, n_274, n_275);
  xor g646 (n_280, n_711, n_276);
  nand g647 (n_712, n_274, n_275);
  nand g648 (n_713, n_276, n_275);
  nand g649 (n_714, n_274, n_276);
  nand g650 (n_301, n_712, n_713, n_714);
  xor g651 (n_715, n_277, n_278);
  xor g652 (n_283, n_715, n_279);
  nand g653 (n_716, n_277, n_278);
  nand g654 (n_717, n_279, n_278);
  nand g655 (n_718, n_277, n_279);
  nand g656 (n_302, n_716, n_717, n_718);
  xor g657 (n_719, n_280, n_281);
  xor g658 (n_285, n_719, n_282);
  nand g659 (n_720, n_280, n_281);
  nand g660 (n_721, n_282, n_281);
  nand g661 (n_722, n_280, n_282);
  nand g662 (n_305, n_720, n_721, n_722);
  xor g663 (n_723, n_283, n_284);
  xor g664 (n_114, n_723, n_285);
  nand g665 (n_724, n_283, n_284);
  nand g666 (n_725, n_285, n_284);
  nand g667 (n_726, n_283, n_285);
  nand g668 (n_92, n_724, n_725, n_726);
  nand g674 (n_308, n_728, n_729, n_730);
  xor g675 (n_731, in_0[8], in_2[7]);
  nand g677 (n_732, in_0[8], in_2[7]);
  nand g680 (n_309, n_732, n_733, n_734);
  xor g682 (n_293, n_735, in_2[10]);
  nand g685 (n_738, in_1[7], in_2[10]);
  nand g686 (n_311, n_736, n_737, n_738);
  xor g687 (n_739, in_2[14], in_1[8]);
  xor g688 (n_295, n_739, in_0[7]);
  nand g689 (n_740, in_2[14], in_1[8]);
  nand g690 (n_741, in_0[7], in_1[8]);
  nand g691 (n_742, in_2[14], in_0[7]);
  nand g692 (n_310, n_740, n_741, n_742);
  xor g693 (n_743, n_288, n_289);
  xor g694 (n_298, n_743, n_290);
  nand g695 (n_744, n_288, n_289);
  nand g696 (n_745, n_290, n_289);
  nand g697 (n_746, n_288, n_290);
  nand g698 (n_316, n_744, n_745, n_746);
  xor g699 (n_747, n_291, n_292);
  xor g700 (n_299, n_747, n_293);
  nand g701 (n_748, n_291, n_292);
  nand g702 (n_749, n_293, n_292);
  nand g703 (n_750, n_291, n_293);
  nand g704 (n_317, n_748, n_749, n_750);
  xor g705 (n_751, n_294, n_295);
  xor g706 (n_300, n_751, n_296);
  nand g707 (n_752, n_294, n_295);
  nand g708 (n_753, n_296, n_295);
  nand g709 (n_754, n_294, n_296);
  nand g710 (n_321, n_752, n_753, n_754);
  xor g711 (n_755, n_297, n_298);
  xor g712 (n_303, n_755, n_299);
  nand g713 (n_756, n_297, n_298);
  nand g714 (n_757, n_299, n_298);
  nand g715 (n_758, n_297, n_299);
  nand g716 (n_322, n_756, n_757, n_758);
  xor g717 (n_759, n_300, n_301);
  xor g718 (n_304, n_759, n_302);
  nand g719 (n_760, n_300, n_301);
  nand g720 (n_761, n_302, n_301);
  nand g721 (n_762, n_300, n_302);
  nand g722 (n_325, n_760, n_761, n_762);
  xor g723 (n_763, n_303, n_304);
  xor g724 (n_113, n_763, n_305);
  nand g725 (n_764, n_303, n_304);
  nand g726 (n_765, n_305, n_304);
  nand g727 (n_766, n_303, n_305);
  nand g728 (n_91, n_764, n_765, n_766);
  nand g734 (n_328, n_768, n_769, n_770);
  xor g735 (n_771, in_0[9], in_2[8]);
  nand g737 (n_772, in_0[9], in_2[8]);
  nand g740 (n_329, n_772, n_773, n_774);
  xor g742 (n_313, n_775, in_2[11]);
  nand g745 (n_778, in_1[8], in_2[11]);
  nand g746 (n_331, n_776, n_777, n_778);
  xor g747 (n_779, in_2[15], in_1[9]);
  xor g748 (n_315, n_779, in_0[8]);
  nand g749 (n_780, in_2[15], in_1[9]);
  nand g750 (n_781, in_0[8], in_1[9]);
  nand g751 (n_782, in_2[15], in_0[8]);
  nand g752 (n_330, n_780, n_781, n_782);
  xor g753 (n_783, n_308, n_309);
  xor g754 (n_318, n_783, n_310);
  nand g755 (n_784, n_308, n_309);
  nand g756 (n_785, n_310, n_309);
  nand g757 (n_786, n_308, n_310);
  nand g758 (n_336, n_784, n_785, n_786);
  xor g759 (n_787, n_311, n_312);
  xor g760 (n_319, n_787, n_313);
  nand g761 (n_788, n_311, n_312);
  nand g762 (n_789, n_313, n_312);
  nand g763 (n_790, n_311, n_313);
  nand g764 (n_337, n_788, n_789, n_790);
  xor g765 (n_791, n_314, n_315);
  xor g766 (n_320, n_791, n_316);
  nand g767 (n_792, n_314, n_315);
  nand g768 (n_793, n_316, n_315);
  nand g769 (n_794, n_314, n_316);
  nand g770 (n_341, n_792, n_793, n_794);
  xor g771 (n_795, n_317, n_318);
  xor g772 (n_323, n_795, n_319);
  nand g773 (n_796, n_317, n_318);
  nand g774 (n_797, n_319, n_318);
  nand g775 (n_798, n_317, n_319);
  nand g776 (n_342, n_796, n_797, n_798);
  xor g777 (n_799, n_320, n_321);
  xor g778 (n_324, n_799, n_322);
  nand g779 (n_800, n_320, n_321);
  nand g780 (n_801, n_322, n_321);
  nand g781 (n_802, n_320, n_322);
  nand g782 (n_345, n_800, n_801, n_802);
  xor g783 (n_803, n_323, n_324);
  xor g784 (n_112, n_803, n_325);
  nand g785 (n_804, n_323, n_324);
  nand g786 (n_805, n_325, n_324);
  nand g787 (n_806, n_323, n_325);
  nand g788 (n_90, n_804, n_805, n_806);
  nand g794 (n_348, n_808, n_809, n_810);
  xor g795 (n_811, in_0[10], in_2[9]);
  nand g797 (n_812, in_0[10], in_2[9]);
  nand g800 (n_349, n_812, n_813, n_814);
  xor g802 (n_333, n_815, in_2[12]);
  nand g805 (n_818, in_1[9], in_2[12]);
  nand g806 (n_351, n_816, n_817, n_818);
  xor g807 (n_819, in_2[16], in_1[10]);
  xor g808 (n_335, n_819, in_0[9]);
  nand g809 (n_820, in_2[16], in_1[10]);
  nand g810 (n_821, in_0[9], in_1[10]);
  nand g811 (n_822, in_2[16], in_0[9]);
  nand g812 (n_350, n_820, n_821, n_822);
  xor g813 (n_823, n_328, n_329);
  xor g814 (n_338, n_823, n_330);
  nand g815 (n_824, n_328, n_329);
  nand g816 (n_825, n_330, n_329);
  nand g817 (n_826, n_328, n_330);
  nand g818 (n_356, n_824, n_825, n_826);
  xor g819 (n_827, n_331, n_332);
  xor g820 (n_339, n_827, n_333);
  nand g821 (n_828, n_331, n_332);
  nand g822 (n_829, n_333, n_332);
  nand g823 (n_830, n_331, n_333);
  nand g824 (n_357, n_828, n_829, n_830);
  xor g825 (n_831, n_334, n_335);
  xor g826 (n_340, n_831, n_336);
  nand g827 (n_832, n_334, n_335);
  nand g828 (n_833, n_336, n_335);
  nand g829 (n_834, n_334, n_336);
  nand g830 (n_361, n_832, n_833, n_834);
  xor g831 (n_835, n_337, n_338);
  xor g832 (n_343, n_835, n_339);
  nand g833 (n_836, n_337, n_338);
  nand g834 (n_837, n_339, n_338);
  nand g835 (n_838, n_337, n_339);
  nand g836 (n_362, n_836, n_837, n_838);
  xor g837 (n_839, n_340, n_341);
  xor g838 (n_344, n_839, n_342);
  nand g839 (n_840, n_340, n_341);
  nand g840 (n_841, n_342, n_341);
  nand g841 (n_842, n_340, n_342);
  nand g842 (n_365, n_840, n_841, n_842);
  xor g843 (n_843, n_343, n_344);
  xor g844 (n_111, n_843, n_345);
  nand g845 (n_844, n_343, n_344);
  nand g846 (n_845, n_345, n_344);
  nand g847 (n_846, n_343, n_345);
  nand g848 (n_89, n_844, n_845, n_846);
  nand g854 (n_368, n_848, n_849, n_850);
  xor g855 (n_851, in_0[11], in_2[10]);
  nand g857 (n_852, in_0[11], in_2[10]);
  nand g860 (n_369, n_852, n_853, n_854);
  xor g862 (n_353, n_855, in_2[13]);
  nand g865 (n_858, in_1[10], in_2[13]);
  nand g866 (n_371, n_856, n_857, n_858);
  xor g867 (n_859, in_2[17], in_1[11]);
  xor g868 (n_355, n_859, in_0[10]);
  nand g869 (n_860, in_2[17], in_1[11]);
  nand g870 (n_861, in_0[10], in_1[11]);
  nand g871 (n_862, in_2[17], in_0[10]);
  nand g872 (n_370, n_860, n_861, n_862);
  xor g873 (n_863, n_348, n_349);
  xor g874 (n_358, n_863, n_350);
  nand g875 (n_864, n_348, n_349);
  nand g876 (n_865, n_350, n_349);
  nand g877 (n_866, n_348, n_350);
  nand g878 (n_376, n_864, n_865, n_866);
  xor g879 (n_867, n_351, n_352);
  xor g880 (n_359, n_867, n_353);
  nand g881 (n_868, n_351, n_352);
  nand g882 (n_869, n_353, n_352);
  nand g883 (n_870, n_351, n_353);
  nand g884 (n_377, n_868, n_869, n_870);
  xor g885 (n_871, n_354, n_355);
  xor g886 (n_360, n_871, n_356);
  nand g887 (n_872, n_354, n_355);
  nand g888 (n_873, n_356, n_355);
  nand g889 (n_874, n_354, n_356);
  nand g890 (n_381, n_872, n_873, n_874);
  xor g891 (n_875, n_357, n_358);
  xor g892 (n_363, n_875, n_359);
  nand g893 (n_876, n_357, n_358);
  nand g894 (n_877, n_359, n_358);
  nand g895 (n_878, n_357, n_359);
  nand g896 (n_382, n_876, n_877, n_878);
  xor g897 (n_879, n_360, n_361);
  xor g898 (n_364, n_879, n_362);
  nand g899 (n_880, n_360, n_361);
  nand g900 (n_881, n_362, n_361);
  nand g901 (n_882, n_360, n_362);
  nand g902 (n_385, n_880, n_881, n_882);
  xor g903 (n_883, n_363, n_364);
  xor g904 (n_110, n_883, n_365);
  nand g905 (n_884, n_363, n_364);
  nand g906 (n_885, n_365, n_364);
  nand g907 (n_886, n_363, n_365);
  nand g908 (n_88, n_884, n_885, n_886);
  nand g914 (n_389, n_888, n_889, n_890);
  xor g915 (n_891, in_0[12], in_2[11]);
  nand g917 (n_892, in_0[12], in_2[11]);
  nand g920 (n_390, n_892, n_893, n_894);
  xor g922 (n_373, n_895, in_2[14]);
  nand g925 (n_898, in_1[11], in_2[14]);
  nand g926 (n_391, n_896, n_897, n_898);
  xor g927 (n_899, in_2[18], in_1[12]);
  xor g928 (n_375, n_899, in_0[11]);
  nand g929 (n_900, in_2[18], in_1[12]);
  nand g930 (n_901, in_0[11], in_1[12]);
  nand g931 (n_902, in_2[18], in_0[11]);
  nand g932 (n_392, n_900, n_901, n_902);
  xor g933 (n_903, n_368, n_369);
  xor g934 (n_378, n_903, n_370);
  nand g935 (n_904, n_368, n_369);
  nand g936 (n_905, n_370, n_369);
  nand g937 (n_906, n_368, n_370);
  nand g938 (n_397, n_904, n_905, n_906);
  xor g939 (n_907, n_371, n_372);
  xor g940 (n_379, n_907, n_373);
  nand g941 (n_908, n_371, n_372);
  nand g942 (n_909, n_373, n_372);
  nand g943 (n_910, n_371, n_373);
  nand g944 (n_399, n_908, n_909, n_910);
  xor g945 (n_911, n_374, n_375);
  xor g946 (n_380, n_911, n_376);
  nand g947 (n_912, n_374, n_375);
  nand g948 (n_913, n_376, n_375);
  nand g949 (n_914, n_374, n_376);
  nand g950 (n_401, n_912, n_913, n_914);
  xor g951 (n_915, n_377, n_378);
  xor g952 (n_383, n_915, n_379);
  nand g953 (n_916, n_377, n_378);
  nand g954 (n_917, n_379, n_378);
  nand g955 (n_918, n_377, n_379);
  nand g956 (n_403, n_916, n_917, n_918);
  xor g957 (n_919, n_380, n_381);
  xor g958 (n_384, n_919, n_382);
  nand g959 (n_920, n_380, n_381);
  nand g960 (n_921, n_382, n_381);
  nand g961 (n_922, n_380, n_382);
  nand g962 (n_406, n_920, n_921, n_922);
  xor g963 (n_923, n_383, n_384);
  xor g964 (n_109, n_923, n_385);
  nand g965 (n_924, n_383, n_384);
  nand g966 (n_925, n_385, n_384);
  nand g967 (n_926, n_383, n_385);
  nand g968 (n_87, n_924, n_925, n_926);
  xor g972 (n_395, n_928, in_2[10]);
  xor g977 (n_933, in_2[19], in_2[15]);
  xor g978 (n_394, n_933, in_0[13]);
  xor g989 (n_943, in_1[12], in_0[12]);
  xor g995 (n_948, n_389, n_390);
  xor g996 (n_398, n_948, n_391);
  xor g1001 (n_953, n_392, n_393);
  xor g1002 (n_400, n_953, n_394);
  xor g1007 (n_958, n_395, n_396);
  xor g1008 (n_402, n_958, n_397);
  xor g1013 (n_963, n_398, n_399);
  xor g1014 (n_404, n_963, n_400);
  xor g1019 (n_968, n_401, n_402);
  xor g1020 (n_405, n_968, n_403);
  xor g1025 (n_973, n_404, n_405);
  xor g1026 (n_108, n_973, n_406);
  nor g1040 (n_993, n_105, n_126);
  nand g1041 (n_988, n_105, n_126);
  nor g1042 (n_989, n_104, n_125);
  nand g1043 (n_990, n_104, n_125);
  nor g1044 (n_999, n_103, n_124);
  nand g1045 (n_994, n_103, n_124);
  nor g1046 (n_995, n_102, n_123);
  nand g1047 (n_996, n_102, n_123);
  nor g1048 (n_1005, n_101, n_122);
  nand g1049 (n_1000, n_101, n_122);
  nor g1050 (n_1001, n_100, n_121);
  nand g1051 (n_1002, n_100, n_121);
  nor g1052 (n_1011, n_99, n_120);
  nand g1053 (n_1006, n_99, n_120);
  nor g1054 (n_1007, n_98, n_119);
  nand g1055 (n_1008, n_98, n_119);
  nor g1056 (n_1017, n_97, n_118);
  nand g1057 (n_1012, n_97, n_118);
  nor g1058 (n_1013, n_96, n_117);
  nand g1059 (n_1014, n_96, n_117);
  nor g1060 (n_1023, n_95, n_116);
  nand g1061 (n_1018, n_95, n_116);
  nor g1062 (n_1019, n_94, n_115);
  nand g1063 (n_1020, n_94, n_115);
  nor g1064 (n_1029, n_93, n_114);
  nand g1065 (n_1024, n_93, n_114);
  nor g1066 (n_1025, n_92, n_113);
  nand g1067 (n_1026, n_92, n_113);
  nor g1068 (n_1035, n_91, n_112);
  nand g1069 (n_1030, n_91, n_112);
  nor g1070 (n_1031, n_90, n_111);
  nand g42 (n_1032, n_90, n_111);
  nor g43 (n_1041, n_89, n_110);
  nand g44 (n_1036, n_89, n_110);
  nor g45 (n_1037, n_88, n_109);
  nand g46 (n_1038, n_88, n_109);
  nand g51 (n_1042, n_986, n_987);
  nor g52 (n_991, n_988, n_989);
  nor g55 (n_1045, n_993, n_989);
  nor g56 (n_997, n_994, n_995);
  nor g59 (n_1051, n_999, n_995);
  nor g60 (n_1003, n_1000, n_1001);
  nor g63 (n_1053, n_1005, n_1001);
  nor g64 (n_1009, n_1006, n_1007);
  nor g67 (n_1061, n_1011, n_1007);
  nor g68 (n_1015, n_1012, n_1013);
  nor g71 (n_1063, n_1017, n_1013);
  nor g72 (n_1021, n_1018, n_1019);
  nor g75 (n_1071, n_1023, n_1019);
  nor g76 (n_1027, n_1024, n_1025);
  nor g79 (n_1073, n_1029, n_1025);
  nor g80 (n_1033, n_1030, n_1031);
  nor g83 (n_1081, n_1035, n_1031);
  nor g84 (n_1039, n_1036, n_1037);
  nor g87 (n_1083, n_1041, n_1037);
  nand g90 (n_1154, n_988, n_1044);
  nand g91 (n_1047, n_1045, n_1042);
  nand g92 (n_1088, n_1046, n_1047);
  nor g93 (n_1049, n_1005, n_1048);
  nand g102 (n_1096, n_1051, n_1053);
  nor g103 (n_1059, n_1017, n_1058);
  nand g112 (n_1103, n_1061, n_1063);
  nor g113 (n_1069, n_1029, n_1068);
  nand g122 (n_1111, n_1071, n_1073);
  nor g123 (n_1079, n_1041, n_1078);
  nand g132 (n_1118, n_1081, n_1083);
  nand g135 (n_1158, n_994, n_1090);
  nand g136 (n_1091, n_1051, n_1088);
  nand g137 (n_1160, n_1048, n_1091);
  nand g140 (n_1163, n_1094, n_1095);
  nand g143 (n_1119, n_1098, n_1099);
  nor g144 (n_1101, n_1023, n_1100);
  nor g147 (n_1129, n_1023, n_1103);
  nor g153 (n_1109, n_1107, n_1100);
  nor g156 (n_1135, n_1103, n_1107);
  nor g157 (n_1113, n_1111, n_1100);
  nor g160 (n_1138, n_1103, n_1111);
  nand g167 (n_1167, n_1006, n_1121);
  nand g168 (n_1122, n_1061, n_1119);
  nand g169 (n_1169, n_1058, n_1122);
  nand g172 (n_1172, n_1125, n_1126);
  nand g175 (n_1175, n_1100, n_1128);
  nand g176 (n_1131, n_1129, n_1119);
  nand g177 (n_1178, n_1130, n_1131);
  nand g178 (n_1134, n_1132, n_1119);
  nand g179 (n_1180, n_1133, n_1134);
  nand g180 (n_1137, n_1135, n_1119);
  nand g181 (n_1183, n_1136, n_1137);
  nand g182 (n_1140, n_1138, n_1119);
  nand g183 (n_1141, n_1139, n_1140);
  nand g1072 (n_1187, n_1030, n_1143);
  nand g1073 (n_1144, n_1081, n_1141);
  nand g1074 (n_1189, n_1078, n_1144);
  nand g1077 (n_1192, n_1147, n_1148);
  nand g1080 (n_1195, n_1116, n_1150);
  xnor g1084 (out_0[2], n_1042, n_1152);
  xnor g1087 (out_0[3], n_1154, n_1155);
  xnor g1089 (out_0[4], n_1088, n_1156);
  xnor g1092 (out_0[5], n_1158, n_1159);
  xnor g1094 (out_0[6], n_1160, n_1161);
  xnor g1097 (out_0[7], n_1163, n_1164);
  xnor g1099 (out_0[8], n_1119, n_1165);
  xnor g1102 (out_0[9], n_1167, n_1168);
  xnor g1104 (out_0[10], n_1169, n_1170);
  xnor g1107 (out_0[11], n_1172, n_1173);
  xnor g1110 (out_0[12], n_1175, n_1176);
  xnor g1113 (out_0[13], n_1178, n_1179);
  xnor g1115 (out_0[14], n_1180, n_1181);
  xnor g1118 (out_0[15], n_1183, n_1184);
  xnor g1120 (out_0[16], n_1141, n_1185);
  xnor g1123 (out_0[17], n_1187, n_1188);
  xnor g1125 (out_0[18], n_1189, n_1190);
  xnor g1128 (out_0[19], n_1192, n_1193);
  xnor g1131 (out_0[20], n_1195, n_1196);
  or g1135 (n_410, wc, in_0[1]);
  not gc (wc, in_2[0]);
  xnor g1136 (n_411, in_0[2], in_2[1]);
  or g1137 (n_412, wc0, in_0[2]);
  not gc0 (wc0, in_2[1]);
  or g1138 (n_413, wc1, in_1[2]);
  not gc1 (wc1, in_2[1]);
  or g1139 (n_414, in_0[2], in_1[2]);
  or g1141 (n_416, wc2, in_0[3]);
  not gc2 (wc2, in_2[2]);
  or g1142 (n_417, wc3, in_1[3]);
  not gc3 (wc3, in_2[2]);
  or g1143 (n_418, in_0[3], in_1[3]);
  xnor g1144 (n_419, in_0[4], in_2[3]);
  or g1145 (n_420, wc4, in_0[4]);
  not gc4 (wc4, in_2[3]);
  or g1146 (n_421, wc5, in_1[0]);
  not gc5 (wc5, in_2[3]);
  or g1147 (n_422, in_0[4], in_1[0]);
  xor g1148 (n_423, in_0[0], in_1[4]);
  or g1149 (n_424, in_0[0], in_1[4]);
  xnor g1150 (n_427, in_1[5], in_2[4]);
  or g1151 (n_428, wc6, in_1[5]);
  not gc6 (wc6, in_2[4]);
  or g1152 (n_429, in_1[5], in_1[1]);
  or g1153 (n_430, wc7, in_1[1]);
  not gc7 (wc7, in_2[4]);
  xnor g1154 (n_431, in_0[1], in_2[0]);
  xnor g1155 (n_439, in_0[6], in_2[1]);
  or g1156 (n_440, wc8, in_0[6]);
  not gc8 (wc8, in_2[1]);
  or g1157 (n_441, wc9, in_1[6]);
  not gc9 (wc9, in_2[1]);
  or g1158 (n_442, in_0[6], in_1[6]);
  xnor g1159 (n_443, in_1[2], in_2[5]);
  or g1160 (n_444, wc10, in_1[2]);
  not gc10 (wc10, in_2[5]);
  or g1161 (n_446, wc11, in_0[2]);
  not gc11 (wc11, in_2[5]);
  xnor g1162 (n_455, in_0[7], in_2[2]);
  or g1163 (n_456, wc12, in_0[7]);
  not gc12 (wc12, in_2[2]);
  or g1164 (n_458, in_0[7], in_0[3]);
  xor g1165 (n_459, in_1[7], in_1[3]);
  or g1166 (n_460, in_1[7], in_1[3]);
  or g1167 (n_461, wc13, in_1[3]);
  not gc13 (wc13, in_1[0]);
  or g1168 (n_462, wc14, in_1[7]);
  not gc14 (wc14, in_1[0]);
  xnor g1169 (n_475, in_0[8], in_2[0]);
  or g1170 (n_476, wc15, in_0[8]);
  not gc15 (wc15, in_2[0]);
  or g1171 (n_477, wc16, in_1[8]);
  not gc16 (wc16, in_2[0]);
  or g1172 (n_478, in_0[8], in_1[8]);
  or g1173 (n_482, wc17, in_0[4]);
  not gc17 (wc17, in_0[0]);
  xnor g1174 (n_483, in_1[4], in_1[1]);
  or g1175 (n_484, wc18, in_1[4]);
  not gc18 (wc18, in_1[1]);
  or g1176 (n_485, wc19, in_1[4]);
  not gc19 (wc19, in_2[7]);
  xnor g1177 (n_503, in_0[9], in_2[1]);
  or g1178 (n_504, wc20, in_0[9]);
  not gc20 (wc20, in_2[1]);
  or g1179 (n_505, wc21, in_1[9]);
  not gc21 (wc21, in_2[1]);
  or g1180 (n_506, in_0[9], in_1[9]);
  or g1182 (n_508, wc22, in_0[5]);
  not gc22 (wc22, in_2[4]);
  or g1183 (n_510, wc23, in_0[5]);
  not gc23 (wc23, in_0[1]);
  xnor g1184 (n_511, in_1[5], in_1[2]);
  or g1185 (n_512, wc24, in_1[5]);
  not gc24 (wc24, in_1[2]);
  or g1186 (n_513, wc25, in_1[5]);
  not gc25 (wc25, in_2[8]);
  xnor g1187 (n_535, in_0[10], in_2[0]);
  or g1188 (n_536, wc26, in_0[10]);
  not gc26 (wc26, in_2[0]);
  or g1189 (n_537, wc27, in_1[6]);
  not gc27 (wc27, in_2[0]);
  or g1190 (n_538, in_0[10], in_1[6]);
  xnor g1191 (n_196, n_539, in_1[10]);
  or g1192 (n_541, wc28, in_1[10]);
  not gc28 (wc28, in_2[2]);
  or g1193 (n_542, in_1[10], wc29);
  not gc29 (wc29, in_0[3]);
  xnor g1194 (n_543, in_0[6], in_1[2]);
  or g1195 (n_544, wc30, in_0[6]);
  not gc30 (wc30, in_1[2]);
  or g1196 (n_545, wc31, in_0[6]);
  not gc31 (wc31, in_2[5]);
  xnor g1197 (n_209, in_0[11], in_2[1]);
  and g1198 (n_228, in_2[1], wc32);
  not gc32 (wc32, in_0[11]);
  xnor g1199 (n_571, in_0[4], in_1[7]);
  or g1200 (n_572, in_1[7], wc33);
  not gc33 (wc33, in_0[4]);
  or g1201 (n_574, wc34, in_1[7]);
  not gc34 (wc34, in_2[3]);
  xnor g1202 (n_575, in_1[11], in_1[3]);
  or g1203 (n_576, wc35, in_1[11]);
  not gc35 (wc35, in_1[3]);
  or g1204 (n_577, wc36, in_0[7]);
  not gc36 (wc36, in_1[3]);
  or g1205 (n_578, in_0[7], in_1[11]);
  xnor g1206 (n_607, in_0[12], in_2[2]);
  or g1207 (n_608, wc37, in_0[12]);
  not gc37 (wc37, in_2[2]);
  or g1208 (n_609, wc38, in_1[8]);
  not gc38 (wc38, in_2[2]);
  or g1209 (n_610, in_0[12], in_1[8]);
  xnor g1210 (n_233, n_611, in_1[12]);
  or g1211 (n_613, wc39, in_1[12]);
  not gc39 (wc39, in_2[4]);
  or g1212 (n_614, in_1[12], wc40);
  not gc40 (wc40, in_0[5]);
  xnor g1213 (n_615, in_0[8], in_1[4]);
  or g1214 (n_616, wc41, in_0[8]);
  not gc41 (wc41, in_1[4]);
  or g1215 (n_617, wc42, in_0[8]);
  not gc42 (wc42, in_2[7]);
  xnor g1216 (n_647, in_0[13], in_2[3]);
  or g1217 (n_648, wc43, in_0[13]);
  not gc43 (wc43, in_2[3]);
  or g1218 (n_649, wc44, in_1[9]);
  not gc44 (wc44, in_2[3]);
  or g1219 (n_650, in_0[13], in_1[9]);
  xnor g1220 (n_252, n_651, in_1[13]);
  or g1221 (n_653, wc45, in_1[13]);
  not gc45 (wc45, in_2[5]);
  or g1222 (n_654, in_1[13], wc46);
  not gc46 (wc46, in_0[6]);
  xnor g1223 (n_655, in_0[9], in_1[5]);
  or g1224 (n_656, wc47, in_0[9]);
  not gc47 (wc47, in_1[5]);
  or g1225 (n_657, wc48, in_0[9]);
  not gc48 (wc48, in_2[8]);
  xnor g1226 (n_687, in_0[14], in_2[4]);
  or g1227 (n_688, wc49, in_0[14]);
  not gc49 (wc49, in_2[4]);
  or g1228 (n_689, wc50, in_1[10]);
  not gc50 (wc50, in_2[4]);
  or g1229 (n_690, in_0[14], in_1[10]);
  xnor g1230 (n_272, n_691, in_1[14]);
  or g1231 (n_693, wc51, in_1[14]);
  not gc51 (wc51, in_2[6]);
  or g1232 (n_694, in_1[14], wc52);
  not gc52 (wc52, in_0[7]);
  xnor g1233 (n_695, in_0[10], in_1[6]);
  or g1234 (n_696, wc53, in_0[10]);
  not gc53 (wc53, in_1[6]);
  or g1235 (n_697, wc54, in_0[10]);
  not gc54 (wc54, in_2[9]);
  xnor g1236 (n_727, in_0[15], in_2[5]);
  or g1237 (n_728, wc55, in_0[15]);
  not gc55 (wc55, in_2[5]);
  or g1238 (n_729, wc56, in_1[11]);
  not gc56 (wc56, in_2[5]);
  or g1239 (n_730, in_0[15], in_1[11]);
  xnor g1240 (n_292, n_731, in_1[15]);
  or g1241 (n_733, wc57, in_1[15]);
  not gc57 (wc57, in_2[7]);
  or g1242 (n_734, in_1[15], wc58);
  not gc58 (wc58, in_0[8]);
  xnor g1243 (n_735, in_0[11], in_1[7]);
  or g1244 (n_736, wc59, in_0[11]);
  not gc59 (wc59, in_1[7]);
  or g1245 (n_737, wc60, in_0[11]);
  not gc60 (wc60, in_2[10]);
  xnor g1246 (n_767, in_0[16], in_2[6]);
  or g1247 (n_768, wc61, in_0[16]);
  not gc61 (wc61, in_2[6]);
  or g1248 (n_769, wc62, in_1[12]);
  not gc62 (wc62, in_2[6]);
  or g1249 (n_770, in_0[16], in_1[12]);
  xnor g1250 (n_312, n_771, in_1[16]);
  or g1251 (n_773, wc63, in_1[16]);
  not gc63 (wc63, in_2[8]);
  or g1252 (n_774, in_1[16], wc64);
  not gc64 (wc64, in_0[9]);
  xnor g1253 (n_775, in_0[12], in_1[8]);
  or g1254 (n_776, wc65, in_0[12]);
  not gc65 (wc65, in_1[8]);
  or g1255 (n_777, wc66, in_0[12]);
  not gc66 (wc66, in_2[11]);
  xnor g1256 (n_807, in_0[17], in_2[7]);
  or g1257 (n_808, wc67, in_0[17]);
  not gc67 (wc67, in_2[7]);
  or g1258 (n_809, wc68, in_1[13]);
  not gc68 (wc68, in_2[7]);
  or g1259 (n_810, in_0[17], in_1[13]);
  xnor g1260 (n_332, n_811, in_1[17]);
  or g1261 (n_813, wc69, in_1[17]);
  not gc69 (wc69, in_2[9]);
  or g1262 (n_814, in_1[17], wc70);
  not gc70 (wc70, in_0[10]);
  xnor g1263 (n_815, in_0[13], in_1[9]);
  or g1264 (n_816, wc71, in_0[13]);
  not gc71 (wc71, in_1[9]);
  or g1265 (n_817, wc72, in_0[13]);
  not gc72 (wc72, in_2[12]);
  xnor g1266 (n_847, in_0[18], in_2[8]);
  or g1267 (n_848, wc73, in_0[18]);
  not gc73 (wc73, in_2[8]);
  or g1268 (n_849, wc74, in_1[14]);
  not gc74 (wc74, in_2[8]);
  or g1269 (n_850, in_0[18], in_1[14]);
  xnor g1270 (n_352, n_851, in_1[18]);
  or g1271 (n_853, wc75, in_1[18]);
  not gc75 (wc75, in_2[10]);
  or g1272 (n_854, in_1[18], wc76);
  not gc76 (wc76, in_0[11]);
  xnor g1273 (n_855, in_0[14], in_1[10]);
  or g1274 (n_856, wc77, in_0[14]);
  not gc77 (wc77, in_1[10]);
  or g1275 (n_857, wc78, in_0[14]);
  not gc78 (wc78, in_2[13]);
  xnor g1276 (n_887, in_0[19], in_2[9]);
  or g1277 (n_888, wc79, in_0[19]);
  not gc79 (wc79, in_2[9]);
  or g1278 (n_889, wc80, in_1[15]);
  not gc80 (wc80, in_2[9]);
  or g1279 (n_890, in_0[19], in_1[15]);
  xnor g1280 (n_372, n_891, in_1[19]);
  or g1281 (n_893, wc81, in_1[19]);
  not gc81 (wc81, in_2[11]);
  or g1282 (n_894, in_1[19], wc82);
  not gc82 (wc82, in_0[12]);
  xnor g1283 (n_895, in_0[15], in_1[11]);
  or g1284 (n_896, wc83, in_0[15]);
  not gc83 (wc83, in_1[11]);
  or g1285 (n_897, wc84, in_0[15]);
  not gc84 (wc84, in_2[14]);
  xnor g1286 (n_928, in_1[16], in_2[12]);
  xnor g1287 (n_938, in_0[16], in_1[13]);
  xnor g1288 (n_396, n_943, in_0[20]);
  or g1289 (n_981, in_0[0], in_1[0]);
  or g1291 (n_105, in_2[0], wc85, wc86);
  not gc86 (wc86, n_410);
  not gc85 (wc85, in_0[1]);
  xnor g1292 (n_126, n_411, in_1[2]);
  xor g1293 (n_125, n_539, in_1[3]);
  xnor g1294 (n_103, n_419, in_1[0]);
  xnor g1295 (n_144, n_427, in_1[1]);
  or g1296 (n_433, in_0[1], wc87);
  not gc87 (wc87, in_0[5]);
  xnor g1297 (n_150, n_439, in_1[6]);
  xnor g1298 (n_151, n_443, in_0[2]);
  xnor g1299 (n_158, n_455, in_0[3]);
  xnor g1300 (n_168, n_475, in_1[8]);
  xnor g1301 (n_180, n_503, in_1[9]);
  xnor g1302 (n_181, n_611, in_0[1]);
  xnor g1303 (n_195, n_535, in_1[6]);
  xnor g1304 (n_215, n_575, in_0[7]);
  xnor g1305 (n_235, n_607, in_1[8]);
  xnor g1306 (n_254, n_647, in_1[9]);
  xnor g1307 (n_274, n_687, in_1[10]);
  xnor g1308 (n_294, n_727, in_1[11]);
  xnor g1309 (n_314, n_767, in_1[12]);
  xnor g1310 (n_334, n_807, in_1[13]);
  xnor g1311 (n_354, n_847, in_1[14]);
  xnor g1312 (n_374, n_887, in_1[15]);
  xnor g1313 (n_393, n_938, in_1[20]);
  xor g1315 (out_0[0], in_0[0], in_1[0]);
  or g1316 (n_425, in_0[0], wc88);
  not gc88 (wc88, n_138);
  or g1317 (n_426, in_1[4], wc89);
  not gc89 (wc89, n_138);
  xnor g1318 (n_447, n_149, in_0[5]);
  or g1319 (n_448, in_0[5], wc90);
  not gc90 (wc90, n_149);
  or g1320 (n_450, in_0[5], wc91);
  not gc91 (wc91, n_150);
  and g1321 (n_983, n_431, in_1[1]);
  or g1322 (n_986, n_431, in_1[1]);
  or g1323 (n_987, n_981, n_983);
  and g1324 (n_1046, wc92, n_990);
  not gc92 (wc92, n_991);
  or g1325 (n_1151, wc93, n_983);
  not gc93 (wc93, n_986);
  or g1326 (n_1152, wc94, n_993);
  not gc94 (wc94, n_988);
  or g1327 (n_1155, wc95, n_989);
  not gc95 (wc95, n_990);
  xor g1328 (out_0[1], n_981, n_1151);
  or g1329 (n_1156, wc96, n_999);
  not gc96 (wc96, n_994);
  and g1330 (n_1048, wc97, n_996);
  not gc97 (wc97, n_997);
  or g1331 (n_1044, wc98, n_993);
  not gc98 (wc98, n_1042);
  or g1332 (n_1159, wc99, n_995);
  not gc99 (wc99, n_996);
  or g1333 (n_1092, wc100, n_1005);
  not gc100 (wc100, n_1051);
  or g1334 (n_1161, wc101, n_1005);
  not gc101 (wc101, n_1000);
  and g1335 (n_1055, wc102, n_1002);
  not gc102 (wc102, n_1003);
  and g1336 (n_1094, wc103, n_1000);
  not gc103 (wc103, n_1049);
  or g1337 (n_1090, wc104, n_999);
  not gc104 (wc104, n_1088);
  or g1338 (n_1164, wc105, n_1001);
  not gc105 (wc105, n_1002);
  and g1339 (n_1056, wc106, n_1053);
  not gc106 (wc106, n_1048);
  or g1340 (n_1095, n_1092, wc107);
  not gc107 (wc107, n_1088);
  or g1341 (n_1165, wc108, n_1011);
  not gc108 (wc108, n_1006);
  and g1342 (n_1058, wc109, n_1008);
  not gc109 (wc109, n_1009);
  and g1343 (n_1098, wc110, n_1055);
  not gc110 (wc110, n_1056);
  or g1344 (n_1123, wc111, n_1017);
  not gc111 (wc111, n_1061);
  or g1345 (n_1099, n_1096, wc112);
  not gc112 (wc112, n_1088);
  or g1346 (n_1168, wc113, n_1007);
  not gc113 (wc113, n_1008);
  or g1347 (n_1170, wc114, n_1017);
  not gc114 (wc114, n_1012);
  and g1348 (n_1115, n_87, n_108);
  or g1349 (n_1117, n_87, n_108);
  and g1350 (n_1065, wc115, n_1014);
  not gc115 (wc115, n_1015);
  and g1351 (n_1068, wc116, n_1020);
  not gc116 (wc116, n_1021);
  and g1352 (n_1075, wc117, n_1026);
  not gc117 (wc117, n_1027);
  and g1353 (n_1078, wc118, n_1032);
  not gc118 (wc118, n_1033);
  and g1354 (n_1085, wc119, n_1038);
  not gc119 (wc119, n_1039);
  and g1355 (n_1125, wc120, n_1012);
  not gc120 (wc120, n_1059);
  or g1356 (n_1107, wc121, n_1029);
  not gc121 (wc121, n_1071);
  or g1357 (n_1145, wc122, n_1041);
  not gc122 (wc122, n_1081);
  or g1358 (n_1121, wc123, n_1011);
  not gc123 (wc123, n_1119);
  or g1359 (n_1126, n_1123, wc124);
  not gc124 (wc124, n_1119);
  or g1360 (n_1173, wc125, n_1013);
  not gc125 (wc125, n_1014);
  or g1361 (n_1176, wc126, n_1023);
  not gc126 (wc126, n_1018);
  or g1362 (n_1179, wc127, n_1019);
  not gc127 (wc127, n_1020);
  or g1363 (n_1181, wc128, n_1029);
  not gc128 (wc128, n_1024);
  or g1364 (n_1184, wc129, n_1025);
  not gc129 (wc129, n_1026);
  or g1365 (n_1185, wc130, n_1035);
  not gc130 (wc130, n_1030);
  or g1366 (n_1188, wc131, n_1031);
  not gc131 (wc131, n_1032);
  or g1367 (n_1190, wc132, n_1041);
  not gc132 (wc132, n_1036);
  or g1368 (n_1193, wc133, n_1037);
  not gc133 (wc133, n_1038);
  and g1369 (n_1066, wc134, n_1063);
  not gc134 (wc134, n_1058);
  and g1370 (n_1076, wc135, n_1073);
  not gc135 (wc135, n_1068);
  and g1371 (n_1086, wc136, n_1083);
  not gc136 (wc136, n_1078);
  and g1372 (n_1132, wc137, n_1071);
  not gc137 (wc137, n_1103);
  or g1373 (n_1196, wc138, n_1115);
  not gc138 (wc138, n_1117);
  and g1374 (n_1100, wc139, n_1065);
  not gc139 (wc139, n_1066);
  and g1375 (n_1108, wc140, n_1024);
  not gc140 (wc140, n_1069);
  and g1376 (n_1112, wc141, n_1075);
  not gc141 (wc141, n_1076);
  and g1377 (n_1147, wc142, n_1036);
  not gc142 (wc142, n_1079);
  and g1378 (n_1116, wc143, n_1085);
  not gc143 (wc143, n_1086);
  or g1379 (n_1128, wc144, n_1103);
  not gc144 (wc144, n_1119);
  and g1380 (n_1105, wc145, n_1071);
  not gc145 (wc145, n_1100);
  and g1381 (n_1130, wc146, n_1018);
  not gc146 (wc146, n_1101);
  and g1382 (n_1133, wc147, n_1068);
  not gc147 (wc147, n_1105);
  and g1383 (n_1136, n_1108, wc148);
  not gc148 (wc148, n_1109);
  and g1384 (n_1139, n_1112, wc149);
  not gc149 (wc149, n_1113);
  or g1385 (n_1143, wc150, n_1035);
  not gc150 (wc150, n_1141);
  or g1386 (n_1148, n_1145, wc151);
  not gc151 (wc151, n_1141);
  or g1387 (n_1150, wc152, n_1118);
  not gc152 (wc152, n_1141);
endmodule

module csa_tree_add_125_31_group_301_GENERIC(in_0, in_1, in_2, out_0);
  input [20:0] in_0;
  input [21:0] in_1, in_2;
  output [20:0] out_0;
  wire [20:0] in_0;
  wire [21:0] in_1, in_2;
  wire [20:0] out_0;
  csa_tree_add_125_31_group_301_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

